-- ID/EX stage registers

-- Accepts control signals and adata from the ID stage.
-- Signals include memory read right, writeback controls, data from Register File
